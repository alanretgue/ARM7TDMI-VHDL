library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Decoder is
    port(
        
    );
end entity Decoder;

architecture Derick of Decoder is
begin

end architecture Derick;